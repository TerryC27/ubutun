module test{

};


endmodule 
