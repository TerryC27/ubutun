module test{

};

always @(posedge clk) begin
	if() begin
		

	end
	else begin

	end
end

endmodule 
