module test{

};

always @(posedge clk) begin
	if() begin

	end
end

endmodule 
