module test{

};

always @(posedge clk) begin
	if() begin
		t= t1;		

	end
	else begin

	end
end

endmodule 
